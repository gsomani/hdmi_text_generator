library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity font_rom is
   port(
      addr: in std_logic_vector(7 downto 0);
      data: out std_logic_vector(7 downto 0)
   );
end font_rom;

architecture arch of font_rom is
   constant ADDR_WIDTH: integer:=8;
   constant DATA_WIDTH: integer:=8;
   type rom_type is array (0 to 2**ADDR_WIDTH-1)
        of std_logic_vector(DATA_WIDTH-1 downto 0);
   -- ROM definition
   constant ROM: rom_type:=(   -- 2^8-by-8
   X"00", -- 0
   X"00", -- 1
   X"7C", -- 2  *****
   X"C6", -- 3 **   **
   X"C6", -- 4 **   **
   X"CE", -- 5 **  ***
   X"DE", -- 6 ** ****
   X"F6", -- 7 **** **
   X"E6", -- 8 ***  **
   X"C6", -- 9 **   **
   X"C6", -- a **   **
   X"7C", -- b  *****
   X"00", -- c
   X"00", -- d
   X"00", -- e
   X"00", -- f
   
   X"00", -- 0
   X"00", -- 1
   X"18", -- 2
   X"38", -- 3
   X"78", -- 4    **
   X"18", -- 5   ***
   X"18", -- 6  ****
   X"18", -- 7    **
   X"18", -- 8    **
   X"18", -- 9    **
   X"18", -- a    **
   X"7E", -- b    **
   X"00", -- c    **
   X"00", -- d  ******
   X"00", -- e
   X"00", -- f 

   X"00", -- 0
   X"00", -- 1
   X"7C", -- 2  *****
   X"C6", -- 3 **   **
   X"06", -- 4      **
   X"0C", -- 5     **
   X"18", -- 6    **
   X"30", -- 7   **
   X"60", -- 8  **
   X"C0", -- 9 **
   X"C6", -- a **   **
   X"FE", -- b *******
   X"00", -- c
   X"00", -- d
   X"00", -- e
   X"00", -- f
   
   X"00", -- 0
   X"00", -- 1
   X"7C", -- 2  *****
   X"C6", -- 3 **   **
   X"06", -- 4      **
   X"06", -- 5      **
   X"3C", -- 6   ****
   X"06", -- 7      **
   X"06", -- 8      **
   X"06", -- 9      **
   X"C6", -- a **   **
   X"7C", -- b  *****
   X"00", -- c
   X"00", -- d
   X"00", -- e
   X"00", -- f
   
   X"00", -- 0
   X"00", -- 1
   X"0C", -- 2     **
   X"1C", -- 3    ***
   X"3C", -- 4   ****
   X"6C", -- 5  ** **
   X"CC", -- 6 **  **
   X"FE", -- 7 *******
   X"0C", -- 8     **
   X"0C", -- 9     **
   X"0C", -- a     **
   X"1E", -- b    ****
   X"00", -- c
   X"00", -- d
   X"00", -- e
   X"00", -- f
   
   X"00", -- 0
   X"00", -- 1
   X"FE", -- 2 *******
   X"C0", -- 3 **
   X"C0", -- 4 **
   X"C0", -- 5 **
   X"FC", -- 6 ******
   X"06", -- 7      **
   X"06", -- 8      **
   X"06", -- 9      **
   X"C6", -- a **   **
   X"7C", -- b  *****
   X"00", -- c
   X"00", -- d
   X"00", -- e
   X"00", -- f
   
   X"00", -- 0
   X"00", -- 1
   X"38", -- 2   ***
   X"60", -- 3  **
   X"C0", -- 4 **
   X"C0", -- 5 **
   X"FC", -- 6 ******
   X"C6", -- 7 **   **
   X"C6", -- 8 **   **
   X"C6", -- 9 **   **
   X"C6", -- a **   **
   X"7C", -- b  *****
   X"00", -- c
   X"00", -- d
   X"00", -- e
   X"00", -- f
   
   X"00", -- 0
   X"00", -- 1
   X"FE", -- 2 *******
   X"C6", -- 3 **   **
   X"06", -- 4      **
   X"06", -- 5      **
   X"0C", -- 6     **
   X"18", -- 7    **
   X"30", -- 8   **
   X"30", -- 9   **
   X"30", -- a   **
   X"30", -- b   **
   X"00", -- c
   X"00", -- d
   X"00", -- e
   X"00", -- f
   
   X"00", -- 0
   X"00", -- 1
   X"7C", -- 2  *****
   X"C6", -- 3 **   **
   X"C6", -- 4 **   **
   X"C6", -- 5 **   **
   X"7C", -- 6  *****
   X"C6", -- 7 **   **
   X"C6", -- 8 **   **
   X"C6", -- 9 **   **
   X"C6", -- a **   **
   X"7C", -- b  *****
   X"00", -- c
   X"00", -- d
   X"00", -- e
   X"00", -- f
   
   X"00", -- 0
   X"00", -- 1
   X"7C", -- 2  *****
   X"C6", -- 3 **   **
   X"C6", -- 4 **   **
   X"C6", -- 5 **   **
   X"7E", -- 6  ******
   X"06", -- 7      **
   X"06", -- 8      **
   X"06", -- 9      **
   X"0C", -- a     **
   X"78", -- b  ****
   X"00", -- c
   X"00", -- d
   X"00", -- e
   X"00", -- f
   
   X"00", -- 0
   X"00", -- 1
   X"10", -- 2    *
   X"38", -- 3   ***
   X"6C", -- 4  ** **
   X"C6", -- 5 **   **
   X"C6", -- 6 **   **
   X"FE", -- 7 *******
   X"C6", -- 8 **   **
   X"C6", -- 9 **   **
   X"C6", -- a **   **
   X"C6", -- b **   **
   X"00", -- c
   X"00", -- d
   X"00", -- e
   X"00", -- f
   
   X"00", -- 0
   X"00", -- 1
   X"FC", -- 2 ******
   X"66", -- 3  **  **
   X"66", -- 4  **  **
   X"66", -- 5  **  **
   X"7C", -- 6  *****
   X"66", -- 7  **  **
   X"66", -- 8  **  **
   X"66", -- 9  **  **
   X"66", -- a  **  **
   X"FC", -- b ******
   X"00", -- c
   X"00", -- d
   X"00", -- e
   X"00", -- f
   
   X"00", -- 0
   X"00", -- 1
   X"3C", -- 2   ****
   X"66", -- 3  **  **
   X"C2", -- 4 **    *
   X"C0", -- 5 **
   X"C0", -- 6 **
   X"C0", -- 7 **
   X"C0", -- 8 **
   X"C2", -- 9 **    *
   X"66", -- a  **  **
   X"3C", -- b   ****
   X"00", -- c
   X"00", -- d
   X"00", -- e
   X"00", -- f
  
   X"00", -- 0
   X"00", -- 1
   X"F8", -- 2 *****
   X"6C", -- 3  ** **
   X"66", -- 4  **  **
   X"66", -- 5  **  **
   X"66", -- 6  **  **
   X"66", -- 7  **  **
   X"66", -- 8  **  **
   X"66", -- 9  **  **
   X"6C", -- a  ** **
   X"F8", -- b *****
   X"00", -- c
   X"00", -- d
   X"00", -- e
   X"00", -- f
  
   X"00", -- 0
   X"00", -- 1
   X"FE", -- 2 *******
   X"66", -- 3  **  **
   X"62", -- 4  **   *
   X"68", -- 5  ** *
   X"78", -- 6  ****
   X"68", -- 7  ** *
   X"60", -- 8  **
   X"62", -- 9  **   *
   X"66", -- a  **  **
   X"FE", -- b *******
   X"00", -- c
   X"00", -- d
   X"00", -- e
   X"00", -- f
   
   X"00", -- 0
   X"00", -- 1
   X"FE", -- 2 *******
   X"66", -- 3  **  **
   X"62", -- 4  **   *
   X"68", -- 5  ** *
   X"78", -- 6  ****
   X"68", -- 7  ** *
   X"60", -- 8  **
   X"60", -- 9  **
   X"60", -- a  **
   X"F0", -- b ****
   X"00", -- c
   X"00", -- d
   X"00", -- e
   X"00" -- f
   );
begin
   data <= ROM(to_integer(unsigned(addr)));
end arch;
